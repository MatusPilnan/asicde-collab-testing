// Go ahead!
